module instruction_memory(input [31:0] in, output [31:0] out);
	reg [31:0] temp;

	always @(in) begin
		case (in)
			32'd0 : temp = 32'b10000000001000000000000000001010;//-- Addi	r1,r0,10
			32'd4 : temp = 32'b00000100010000000000100000000000;//-- Add 	r2,r0,r1
			32'd8 : temp = 32'b00001100011000000000100000000000;//-- sub	r3,r0,r1
			32'd12 : temp = 32'b00010100100000100001100000000000;//-- And	r4,r2,r3
			32'd16 : temp = 32'b10000100101000000000001000110100;//-- Subi	r5,r0,564
			32'd20 : temp = 32'b00011000101001010001100000000000;//-- or	r5,r5,r3
			32'd24 : temp = 32'b00011100110001010000000000000000;//-- nor 	r6,r5,r0
			32'd28 : temp = 32'b00100000000001010000100000000000;//-- xor	r0,r5,r1
			32'd32 : temp = 32'b00100000111001010000000000000000;//-- xor	r7,r5,r0
			32'd36 : temp = 32'b00100100111001000001000000000000;//-- sla	r7,r4,r2
			32'd40 : temp = 32'b00101001000000110001000000000000;//-- sll	r8,r3,r2
			32'd44 : temp = 32'b00101101001001100001000000000000;//-- sra	r9,r6,r2
			32'd48 : temp = 32'b00110001010001100001000000000000;//-- srl	r10,r6,r2
			32'd52 : temp = 32'b10000000001000000000010000000000;//-- Addi 	r1,r0,1024
			32'd56 : temp = 32'b10010100010000010000000000000000;//-- st	r2,r1,0
			32'd60 : temp = 32'b10010001011000010000000000000000;//-- ld	r11,r1,0
			32'd64 : temp = 32'b10010100011000010000000000000100;//-- st	r3,r1,4
			32'd68 : temp = 32'b10010100100000010000000000001000;//-- st	r4,r1,8
			32'd72 : temp = 32'b10010100101000010000000000001100;//-- st	r5,r1,12
			32'd76 : temp = 32'b10010100110000010000000000010000;//-- st	r6,r1,16
			32'd80 : temp = 32'b10010100111000010000000000010100;//-- st	r7,r1,20
			32'd84 : temp = 32'b10010101000000010000000000011000;//-- st	r8,r1,24
			32'd88 : temp = 32'b10010101001000010000000000011100;//-- st	r9,r1,28
			32'd92 : temp = 32'b10010101010000010000000000100000;//-- st	r10,r1,32
			32'd96 : temp = 32'b10010101011000010000000000100100;//-- st	r11,r1,36
			32'd100 : temp = 32'b10000000001000000000000000000011;//-- Addi 	r1,r0,3
			32'd104 : temp = 32'b10000000100000000000010000000000;//-- Addi	r4,r0,1024
			32'd108 : temp = 32'b10000000010000000000000000000000;//-- Addi 	r2,r0,0
			32'd112 : temp = 32'b10000000011000000000000000000001;//-- Addi 	r3,r0,1
			32'd116 : temp = 32'b10000001001000000000000000000010;//-- Addi 	r9,r0,2
			32'd120 : temp = 32'b00101001000000110100100000000000;//-- sll	r8,r3,r9
			32'd124 : temp = 32'b00000101000001000100000000000000;//-- Add 	r8,r4,r8
			32'd128 : temp = 32'b10010000101010000000000000000000;//-- ld	r5,r8,0
			32'd132 : temp = 32'b10010000110010001111111111111100;//-- ld	r6,r8,-4
			32'd136 : temp = 32'b00001101001001010011000000000000;//-- sub 	r9,r5,r6
			32'd140 : temp = 32'b10000001010000001000000000000000;//-- Addi 	r10,r0,0x8000
			32'd144 : temp = 32'b10000001011000000000000000010000;//-- Addi	r11,r0,16
			32'd148 : temp = 32'b00101001010010100101100000000000;//-- sll	r10,r10,r11
			32'd152 : temp = 32'b00010101001010010101000000000000;//-- And 	r9,r9,r10
			32'd156 : temp = 32'b10100000000010010000000000000010;//-- Bez	r9,2 -> 8
			32'd160 : temp = 32'b10010100101010001111111111111100;//-- st	r5,r8,-4
			32'd164 : temp = 32'b10010100110010000000000000000000;//-- st	r6,r8,0
			32'd168 : temp = 32'b10000000011000110000000000000001;//-- Addi 	r3,r3,1
			32'd172 : temp = 32'b10100100011000011111111111110001;//-- BNE	r3,r1,-15 -> -42
			32'd176 : temp = 32'b10000000010000100000000000000001;//-- Addi 	r2,r2,1
			32'd180 : temp = 32'b10100100010000011111111111101110;//-- BNE	r2,r1,-18 -> -51
			32'd184 : temp = 32'b10000000001000000000010000000000;//-- Addi 	r1,r0,1024
			32'd188 : temp = 32'b10010000010000010000000000000000;//-- ld	r2,r1,0
			32'd192 : temp = 32'b10010000011000010000000000000100;//-- ld	r3,r1,4
			32'd196 : temp = 32'b10010000100000010000000000001000;//-- ld	r4,r1,8
			32'd200 : temp = 32'b10010000101000010000000000001100;//-- ld	r5,r1,12
			32'd204 : temp = 32'b10010000110000010000000000010000;//-- ld	r6,r1,16
			32'd208 : temp = 32'b10010000111000010000000000010100;//-- ld	r7,r1,20
			32'd212 : temp = 32'b10010001000000010000000000011000;//-- ld	r8,r1,24
			32'd216 : temp = 32'b10010001001000010000000000011100;//-- ld	r9,r1,28
			32'd220 : temp = 32'b10010001010000010000000000100000;//-- ld	r10,r1,32
			32'd224 : temp = 32'b10010001011000010000000000100100;//-- ld	r11,r1,36
			32'd228 : temp = 32'b10101000000000001111111111111100;//-- JMP 	-4
		endcase
	end

	assign out = temp;
endmodule